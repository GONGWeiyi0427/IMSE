
* Value of the capacitance as a function of x for a capacitive transducer 
* of selectable type
* Input: the displacement (x)
* output : the voltage numerically equal to the value of a capacitance

* Dimension parameters (not used for all types of transducers, see the type parameter definition for the meaning): 
* S, d0, l0, w 
* grad : the direction of the x axis. Can take only two values, 1 and -1.
* If grad is 1: the capacitance increases with x
* If grad is 0: the capacitance decreases as x increases 
* grad parameters is not used for symetric transducers where the function C(x) is pair


* type: the type of the transducer. 
* type=1: gap closing, relevant parameters 
*       -initial gap d0
*       -transducer area S
*       -grad 

* type=2: area overlap, relevant parameters 
*       -gap d0
*       -Initial overlapping length l0
*       -Number of parallel capacitors N
*       -width of the structure in the direction normal to the motion w
*       -grad 

* type=3: Symetrical gap closing, relevant parameters 
*       -initial gap d0
*       -transducer area S

* Default values of all parameters are zero: the user **must** 
* explicitely defind the parameters relevant for the used type

.subckt varcap x capa d0=0 S=0 w=0 l0=0 grad=0 type=0
Bcapa capa 0 v={ (type==1? {8.85e-12*S/(d0-grad*v(x))}:
+                (type==2? {8.85e-12*w*N*(l0+grad*v(x))/d0}}:
+                (type==3? {8.85e-12*S*2*d0/(d0**2-v(x)**2)}:0
+                )))}
.ends

** Integrator : out = integral (in)  
** Parameter : k is the integrator gain, 1 by default
.subckt integrator in out k=1 
** The integrator is implemented with a 1 Farad capacitor
** and a voltage controled current source
*Voltage controled current source
G1 0 out1 in 0 1 
C  out1 0 {1/k} 
** We copy the output voltage with a buffer (a voltage follower)
E1 out 0 out1 0 1
.ends

** Derivator : out = deriv (in)  
.subckt derivator in out k=1 
** The derivator is implemented with a 1 Farad capacitor
** and a current controled voltage source

** Copy of the input 
E1 copy_in 0 in 0 1
C copy_in a1 {k} 
Vampermeter a1 0 0
*Current controled voltage source
H1 out 0 Vampermeter 1 

** An alternative way to implement a derivator: with using an integrator
** and an ideal operational amplifier
*Xinteg out copy_in integrator
*E1 out 0 in copy_in 1e8 

.ends

* This subcircuit models a capacitive transducer 
* x (input): the node whose voltage equals the displacement of the mobile electrode
* f (output): the node whose the voltage equals the force generated by the transducer
* cp, cn : the electrical terminals of a dipole representing the variable capacitor

* the parameters: the same as for the subcircuit capvar 
.subckt transducer x f cp cn capax d0=0 S=0 w=0 l0=0 grad=0 type=0
** internal parameter : variation for calculation of the gradient 
.param dx=1e-8

Xcapax x capax varcap d0={d0} S={S} w={w} l0={l0} grad={grad} type={type}

* Definition of the x + delta x for the space gradient calculation
Vdx xpdx x dx 
* Definition of the value of the transducer capacitor as a function
* of x+ delta x
Xcapaxpdx xpdx capaxpdx varcap d0={d0} S={S} w={w} l0={l0} grad={grad} type={type}

** Calculation of the transducer force
Bforce f 0  v={0.5*V(cp, cn)*V(cp, cn)*(V(capaxpdx)-V(capax))/dx}

** Definition of the transducer charge
Bcharge charge 0 v={v(capax)*v(cp, cn)}
** Calcul du courant du trasnducteur
Xcurrent charge vcurrent derivator 

** Generateur de courant du transducteur
GIcvar cp cn vcurrent 0  1
.ends


** Additionneur à deux entrées  
.subckt adder2 in1 in2 out 
E1 out out1 in1 0 1
E2 out1 0 in2 0 1
.ends

** Additionneur à trois entrées  
.subckt adder3 in1 in2 in3 out 
E1 out out1 in1 0 1
E2 out1 out2 in2 0 1
E3 out2 0 in3 0 1
.ends

** Additionneur à quatre entrées  
.subckt adder4 in1 in2 in3 in4 out 
E1 out out1 in1 0 1
E2 out1 out2 in2 0 1
E3 out2 out3 in3 0 1
E4 out3 0 in4 0 1
.ends


** Résonateur mécanique
.subckt resonator ext_force transd_force displacement  k=0 mass=0 mu=0 

** On modélise l'équation de Newton
** a ==> v ==> x (double intégration)
Xint1 a v integrator
Xint2 v displacement integrator

** on multiplie x par -k
E1 kx 0 displacement 0 {-k} 

** on multiplie v par -mu 
E2 muv 0 v 0 {-mu}

** On additionne toutes les  forces
Xadd4 kx muv ext_force transd_force sum_f adder4

** et on boucle la boucle
E3 a 0 sum_f 0 {1/mass} 
.ends

** Modèle des stoppeurs 
.subckt stopper displacement force dstop=70e-6 kst=1e6 must=1
Xderiv displacement v derivator  
Bforce force 0 v=(abs(V(displacement))<dstop ? {0}: {-kst*(abs(v(displacement))-dstop)*sgn(v(displacement))-must*v(v)})
.ends



